library verilog;
use verilog.vl_types.all;
entity g07_testbed_diagram_vlg_vec_tst is
end g07_testbed_diagram_vlg_vec_tst;
