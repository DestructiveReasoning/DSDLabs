$date
  Mon Mar 27 22:14:27 2017
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$var reg 1 ! clock $end
$var reg 1 " finished $end
$var reg 1 # enable $end
$var reg 1 $ reset $end
$var reg 1 % full $end
$var reg 1 & empty $end
$var reg 2 ' mode[1:0] $end
$var reg 6 ( addr[5:0] $end
$var reg 6 ) num[5:0] $end
$var reg 6 * data[5:0] $end
$var reg 6 + value[5:0] $end
$scope module bjt $end
$var reg 1 , clock $end
$var reg 1 - enable $end
$var reg 1 . reset $end
$var reg 2 / mode[1:0] $end
$var reg 6 0 addr[5:0] $end
$var reg 6 1 data[5:0] $end
$var reg 1 2 full $end
$var reg 1 3 empty $end
$var reg 6 4 num[5:0] $end
$var reg 6 5 value[5:0] $end
$var reg 312 6 memory[311:0] $end
$var reg 1 7 t_full $end
$var reg 1 8 t_empty $end
$var integer 32 9 t_num $end
$upscope $end
$enddefinitions $end
#0
1!
0"
0#
0$
0%
1&
b00 '
b011000 (
b000000 )
b101010 *
b000000 +
1,
0-
0.
b00 /
b011000 0
b101010 1
02
13
b000000 4
b000000 5
b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 6
07
18
b0 9
#10000000
0!
0,
#20000000
1!
1,
#30000000
0!
0,
#40000000
1!
b10 '
1,
b10 /
#50000000
0!
0,
#58000000
1#
1-
#60000000
1!
1%
0&
b110100 )
b011000 +
1,
12
03
b110100 4
b011000 5
b110011110010110001110000101111101110101101101100101011101010101001101000100111100110100101100100100011100010100001100000011111011110011101011100011011011010011001011000010111010110010101010100010011010010010001010000001111001110001101001100001011001010001001001000000111000110000101000100000011000010000001000000 6
17
08
b110100 9
#70000000
0!
0,
#80000000
1!
b011001 (
b011001 +
1,
b011001 0
b011001 5
#90000000
0!
0,
#98000000
b01 '
b01 /
#100000000
1!
1,
#110000000
0!
0,
#118000000
b11 '
b11 /
#120000000
1!
0%
b110011 )
b011010 +
1,
02
b110011 4
b011010 5
b000000110011110010110001110000101111101110101101101100101011101010101001101000100111100110100101100100100011100010100001100000011111011110011101011100011011011010011000010111010110010101010100010011010010010001010000001111001110001101001100001011001010001001001000000111000110000101000100000011000010000001000000 6
07
b110011 9
#130000000
0!
0,
#138000000
b00 '
b011010 (
b011011 +
b00 /
b011010 0
b011011 5
#140000000
1!
1,
#150000000
0!
0,
#158000000
b011000 (
b011000 +
b011000 0
b011000 5
#160000000
1!
1,
#170000000
0!
0,
#178000000
b01 '
b01 /
#180000000
1!
1%
b110100 )
b010111 +
1,
12
b110100 4
b010111 5
b110011110010110001110000101111101110101101101100101011101010101001101000100111100110100101100100100011100010100001100000011111011110011101011100011011011010011000010111010110010101010100010011010010010001010000001111001110001101001100001011001010001001001000000111000110000101000100000011000010000001000000101010 6
17
b110100 9
#190000000
0!
0,
#198000000
b00 '
b000000 (
b101010 +
b00 /
b000000 0
b101010 5
#200000000
1!
1,
#210000000
0!
0,
#218000000
b11 '
b11 /
#220000000
1!
0%
b110011 )
b000000 +
1,
02
b110011 4
b000000 5
b000000110011110010110001110000101111101110101101101100101011101010101001101000100111100110100101100100100011100010100001100000011111011110011101011100011011011010011000010111010110010101010100010011010010010001010000001111001110001101001100001011001010001001001000000111000110000101000100000011000010000001000000 6
07
b110011 9
#230000000
0!
0,
#238000000
b00 '
b00 /
#240000000
1!
1,
#250000000
0!
0,
#258000000
b11 '
b110011 (
b11 /
b110011 0
#260000000
1!
b110010 )
1,
b110010 4
b110010 9
#270000000
0!
0,
#278000000
b00 '
b00 /
#280000000
1!
1,
#290000000
0!
0,
#298000000
b110010 (
b110011 +
b110010 0
b110011 5
#300000000
1!
1,
#301000000
1$
1&
b000000 )
b000000 +
1.
13
b000000 4
b000000 5
b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 6
18
b0 9
#303000000
0$
0.
#310000000
0!
0,
#318000000
b11 '
b111111 (
b11 /
b111111 0
#320000000
1!
1,
#330000000
0!
0,
#338000000
1"
