$date
  Thu Mar 30 16:02:33 2017
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$var reg 1 ! turn $end
$var reg 1 " cnt_lt_num $end
$var reg 1 # valid $end
$var reg 1 $ reset $end
$var reg 1 % stack_enable $end
$var reg 1 & cnt_reg_enable $end
$var reg 1 ' cnt_reset $end
$var reg 1 ( done $end
$var reg 1 ) clock $end
$var reg 1 * finished $end
$var reg 2 + stack_mode[1:0] $end
$scope module fsm $end
$var reg 1 , turn $end
$var reg 1 - cnt_lt_num $end
$var reg 1 . valid $end
$var reg 1 / clock $end
$var reg 1 0 reset $end
$var reg 1 1 stack_enable $end
$var reg 2 2 stack_mode[1:0] $end
$var reg 1 3 cnt_reg_enable $end
$var reg 1 4 cnt_reset $end
$var reg 1 5 done $end
$comment state is not handled $end
$upscope $end
$enddefinitions $end
#0
0!
1"
0#
0$
0%
0&
1'
0(
1)
0*
b00 +
0,
1-
0.
1/
00
01
b00 2
03
14
05
#10000000
0)
0/
#18000000
1!
1,
#20000000
1&
0'
1)
1/
13
04
#30000000
0)
0/
#38000000
1#
1.
#40000000
1%
0&
1(
1)
b11 +
1/
11
b11 2
03
15
#50000000
0)
0/
#58000000
0!
0#
0,
0.
#60000000
0%
1'
0(
1)
b00 +
1/
01
b00 2
14
05
#70000000
0)
0/
#78000000
1!
1,
#80000000
1&
0'
1)
1/
13
04
#90000000
0)
0/
#98000000
0"
0-
#100000000
1%
1)
b01 +
1/
11
b01 2
#110000000
0)
0/
#120000000
1)
1/
#130000000
0)
0/
#138000000
1"
1#
1-
1.
#140000000
0&
1(
1)
b11 +
1/
b11 2
03
15
#150000000
0)
0/
#160000000
0%
1'
0(
1)
b00 +
1/
01
b00 2
14
05
#170000000
0)
0/
#180000000
1&
0'
1)
1/
13
04
#185000000
1$
0&
1'
10
03
14
#187000000
0!
0$
0,
00
#190000000
0)
0/
#198000000
1*
