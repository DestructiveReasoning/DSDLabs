-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.0.0 Build 156 04/24/2013 SJ Web Edition"
-- CREATED		"Thu Feb  2 16:13:02 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY g07_adder IS 
	PORT
	(
		Sub :  IN  STD_LOGIC;
		A :  IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		B :  IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		S :  OUT  STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END g07_adder;

ARCHITECTURE bdf_type OF g07_adder IS 

SIGNAL	S_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(9 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_86 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_87 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_88 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_89 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_90 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_91 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_92 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_93 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_94 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_95 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_96 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_97 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_98 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_99 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_100 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_101 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_102 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_103 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_104 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;


BEGIN 



S_ALTERA_SYNTHESIZED(6) <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_78;


S_ALTERA_SYNTHESIZED(7) <= SYNTHESIZED_WIRE_2 AND SYNTHESIZED_WIRE_78;


S_ALTERA_SYNTHESIZED(8) <= SYNTHESIZED_WIRE_4 AND SYNTHESIZED_WIRE_78;


S_ALTERA_SYNTHESIZED(9) <= SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_78;


SYNTHESIZED_WIRE_80 <= A(0) XOR SYNTHESIZED_WIRE_79;


S_ALTERA_SYNTHESIZED(0) <= Sub XOR SYNTHESIZED_WIRE_80;


SYNTHESIZED_WIRE_83 <= A(2) XOR SYNTHESIZED_WIRE_81;


S_ALTERA_SYNTHESIZED(2) <= SYNTHESIZED_WIRE_82 XOR SYNTHESIZED_WIRE_83;


SYNTHESIZED_WIRE_16 <= A(2) AND SYNTHESIZED_WIRE_81;


SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_82 AND SYNTHESIZED_WIRE_83;


SYNTHESIZED_WIRE_85 <= SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17;


SYNTHESIZED_WIRE_86 <= A(3) XOR SYNTHESIZED_WIRE_84;


S_ALTERA_SYNTHESIZED(3) <= SYNTHESIZED_WIRE_85 XOR SYNTHESIZED_WIRE_86;


SYNTHESIZED_WIRE_24 <= A(3) AND SYNTHESIZED_WIRE_84;


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_85 AND SYNTHESIZED_WIRE_86;


SYNTHESIZED_WIRE_88 <= SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25;


SYNTHESIZED_WIRE_50 <= A(0) AND SYNTHESIZED_WIRE_79;


SYNTHESIZED_WIRE_89 <= A(4) XOR SYNTHESIZED_WIRE_87;


S_ALTERA_SYNTHESIZED(4) <= SYNTHESIZED_WIRE_88 XOR SYNTHESIZED_WIRE_89;


SYNTHESIZED_WIRE_33 <= A(4) AND SYNTHESIZED_WIRE_87;


SYNTHESIZED_WIRE_34 <= SYNTHESIZED_WIRE_88 AND SYNTHESIZED_WIRE_89;


SYNTHESIZED_WIRE_91 <= SYNTHESIZED_WIRE_33 OR SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_92 <= A(5) XOR SYNTHESIZED_WIRE_90;


S_ALTERA_SYNTHESIZED(5) <= SYNTHESIZED_WIRE_91 XOR SYNTHESIZED_WIRE_92;


SYNTHESIZED_WIRE_41 <= A(5) AND SYNTHESIZED_WIRE_90;


SYNTHESIZED_WIRE_42 <= SYNTHESIZED_WIRE_91 AND SYNTHESIZED_WIRE_92;


SYNTHESIZED_WIRE_94 <= SYNTHESIZED_WIRE_41 OR SYNTHESIZED_WIRE_42;


SYNTHESIZED_WIRE_51 <= Sub AND SYNTHESIZED_WIRE_80;


SYNTHESIZED_WIRE_95 <= A(6) XOR SYNTHESIZED_WIRE_93;


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_94 XOR SYNTHESIZED_WIRE_95;


SYNTHESIZED_WIRE_79 <= B(0) XOR Sub;


SYNTHESIZED_WIRE_102 <= B(1) XOR Sub;


SYNTHESIZED_WIRE_81 <= B(2) XOR Sub;


SYNTHESIZED_WIRE_84 <= B(3) XOR Sub;


SYNTHESIZED_WIRE_87 <= B(4) XOR Sub;


SYNTHESIZED_WIRE_90 <= B(5) XOR Sub;


SYNTHESIZED_WIRE_52 <= A(6) AND SYNTHESIZED_WIRE_93;


SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_94 AND SYNTHESIZED_WIRE_95;


SYNTHESIZED_WIRE_103 <= SYNTHESIZED_WIRE_50 OR SYNTHESIZED_WIRE_51;


SYNTHESIZED_WIRE_97 <= SYNTHESIZED_WIRE_52 OR SYNTHESIZED_WIRE_53;


SYNTHESIZED_WIRE_93 <= B(6) XOR Sub;


SYNTHESIZED_WIRE_98 <= A(7) XOR SYNTHESIZED_WIRE_96;


SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_97 XOR SYNTHESIZED_WIRE_98;


SYNTHESIZED_WIRE_74 <= A(7) AND SYNTHESIZED_WIRE_96;


SYNTHESIZED_WIRE_75 <= SYNTHESIZED_WIRE_97 AND SYNTHESIZED_WIRE_98;


SYNTHESIZED_WIRE_101 <= A(8) XOR SYNTHESIZED_WIRE_99;


SYNTHESIZED_WIRE_96 <= B(7) XOR Sub;


SYNTHESIZED_WIRE_78 <= NOT(Sub);



SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_100 XOR SYNTHESIZED_WIRE_101;


SYNTHESIZED_WIRE_104 <= A(1) XOR SYNTHESIZED_WIRE_102;


SYNTHESIZED_WIRE_76 <= A(8) AND SYNTHESIZED_WIRE_99;


SYNTHESIZED_WIRE_77 <= SYNTHESIZED_WIRE_100 AND SYNTHESIZED_WIRE_101;


SYNTHESIZED_WIRE_99 <= B(8) XOR Sub;


S_ALTERA_SYNTHESIZED(1) <= SYNTHESIZED_WIRE_103 XOR SYNTHESIZED_WIRE_104;


SYNTHESIZED_WIRE_72 <= A(1) AND SYNTHESIZED_WIRE_102;


SYNTHESIZED_WIRE_73 <= SYNTHESIZED_WIRE_103 AND SYNTHESIZED_WIRE_104;


SYNTHESIZED_WIRE_82 <= SYNTHESIZED_WIRE_72 OR SYNTHESIZED_WIRE_73;


SYNTHESIZED_WIRE_100 <= SYNTHESIZED_WIRE_74 OR SYNTHESIZED_WIRE_75;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_76 OR SYNTHESIZED_WIRE_77;

S <= S_ALTERA_SYNTHESIZED;

END bdf_type;