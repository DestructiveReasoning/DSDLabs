library verilog;
use verilog.vl_types.all;
entity g07_debounder_vlg_check_tst is
    port(
        PULSE           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g07_debounder_vlg_check_tst;
